/* This is a starting comment */
module Test;
    // This is an inline comment
    wire x; //It starts here, too
endmodule
/* This is an ending comment */


