module First (x);
    input x;
    CSA csa1_0_10(x);
    CSA csa2_10_0(1'b0);
endmodule

module Second (y, z);
    input y;
    output z;

    CSA CSA_10_0(x);
    CSA CSA_80_0(x);
    CSA CSA_160_0(x);
endmodule

module CSA(item);
    input item;

    // Do nothing! Woo!
endmodule

module Third;
    wire [7:0] x;
    wire [3:0] y;
    and2 a00(x[0], x[1], y[0]);
    and2 a01(x[2], x[3], y[1]);
    and2 a02(x[4], x[5], y[2]);
    and2 a03(x[6], x[7], y[3]);
endmodule

module and2(x0, x1, y);
    input x0;
    input x1;
    output y;
endmodule
