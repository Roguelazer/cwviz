module Hello (input x, output [31:0] y);
    // comament
    CSA CSA_0_3(x[1], y[2], z);
endmodule
