//../verilog/arrayFlat/mult_arrayFlat_16_16.v
//this is an automatically generated unsigned array multiplier that is MbyN bits
//It was created by multGenFlat.pl
module multiplier(//An Unsigned M by N Array multiplier
    input   [15:0] x,
    input   [15:0] y,
    output  [31:0] p);

    wire    ip0[0:14];
    wire    ip1[0:14];
    wire    ip2[0:14];
    wire    ip3[0:14];
    wire    ip4[0:14];
    wire    ip5[0:14];
    wire    ip6[0:14];
    wire    ip7[0:14];
    wire    ip8[0:14];
    wire    ip9[0:14];
    wire    ip10[0:14];
    wire    ip11[0:14];
    wire    ip12[0:14];
    wire    ip13[0:14];
    wire    ip14[0:14];
    wire    ip15[0:14];
    wire    c0[0:15];
    wire    c1[0:15];
    wire    c2[0:15];
    wire    c3[0:15];
    wire    c4[0:15];
    wire    c5[0:15];
    wire    c6[0:15];
    wire    c7[0:15];
    wire    c8[0:15];
    wire    c9[0:15];
    wire    c10[0:15];
    wire    c11[0:15];
    wire    c12[0:15];
    wire    c13[0:15];
    wire    c14[0:15];
    wire    c15[0:15];
    wire    c16[0:15];

    CSA     CSA_0_0(c0[0],p  [0],1'b0  ,1'b0 ,x[0],y[0]);
    CSA     CSA_80_0(c0[1],ip0[0],1'b0  ,1'b0 ,x[1],y[0]);
    CSA     CSA_160_0(c0[2],ip0[1],1'b0  ,1'b0 ,x[2],y[0]);
    CSA     CSA_240_0(c0[3],ip0[2],1'b0  ,1'b0 ,x[3],y[0]);
    CSA     CSA_320_0(c0[4],ip0[3],1'b0  ,1'b0 ,x[4],y[0]);
    CSA     CSA_400_0(c0[5],ip0[4],1'b0  ,1'b0 ,x[5],y[0]);
    CSA     CSA_480_0(c0[6],ip0[5],1'b0  ,1'b0 ,x[6],y[0]);
    CSA     CSA_560_0(c0[7],ip0[6],1'b0  ,1'b0 ,x[7],y[0]);
    CSA     CSA_640_0(c0[8],ip0[7],1'b0  ,1'b0 ,x[8],y[0]);
    CSA     CSA_720_0(c0[9],ip0[8],1'b0  ,1'b0 ,x[9],y[0]);
    CSA     CSA_800_0(c0[10],ip0[9],1'b0  ,1'b0 ,x[10],y[0]);
    CSA     CSA_880_0(c0[11],ip0[10],1'b0  ,1'b0 ,x[11],y[0]);
    CSA     CSA_960_0(c0[12],ip0[11],1'b0  ,1'b0 ,x[12],y[0]);
    CSA     CSA_1040_0(c0[13],ip0[12],1'b0  ,1'b0 ,x[13],y[0]);
    CSA     CSA_1120_0(c0[14],ip0[13],1'b0  ,1'b0 ,x[14],y[0]);
    CSA     CSA_1200_0(c0[15],ip0[14],1'b0  ,1'b0 ,x[15],y[0]);
    CSA     CSA_0_168(c1[0],p  [1],ip0[0],c0[0],x[0],y[1]);
    CSA     CSA_80_168(c1[1],ip1[0],ip0[1],c0[1],x[1],y[1]);
    CSA     CSA_160_168(c1[2],ip1[1],ip0[2],c0[2],x[2],y[1]);
    CSA     CSA_240_168(c1[3],ip1[2],ip0[3],c0[3],x[3],y[1]);
    CSA     CSA_320_168(c1[4],ip1[3],ip0[4],c0[4],x[4],y[1]);
    CSA     CSA_400_168(c1[5],ip1[4],ip0[5],c0[5],x[5],y[1]);
    CSA     CSA_480_168(c1[6],ip1[5],ip0[6],c0[6],x[6],y[1]);
    CSA     CSA_560_168(c1[7],ip1[6],ip0[7],c0[7],x[7],y[1]);
    CSA     CSA_640_168(c1[8],ip1[7],ip0[8],c0[8],x[8],y[1]);
    CSA     CSA_720_168(c1[9],ip1[8],ip0[9],c0[9],x[9],y[1]);
    CSA     CSA_800_168(c1[10],ip1[9],ip0[10],c0[10],x[10],y[1]);
    CSA     CSA_880_168(c1[11],ip1[10],ip0[11],c0[11],x[11],y[1]);
    CSA     CSA_960_168(c1[12],ip1[11],ip0[12],c0[12],x[12],y[1]);
    CSA     CSA_1040_168(c1[13],ip1[12],ip0[13],c0[13],x[13],y[1]);
    CSA     CSA_1120_168(c1[14],ip1[13],ip0[14],c0[14],x[14],y[1]);
    CSA     CSA_1200_168(c1[15],ip1[14],1'b0  ,c0[15],x[15],y[1]);
    CSA     CSA_0_336(c2[0],p  [2],ip1[0],c1[0],x[0],y[2]);
    CSA     CSA_80_336(c2[1],ip2[0],ip1[1],c1[1],x[1],y[2]);
    CSA     CSA_160_336(c2[2],ip2[1],ip1[2],c1[2],x[2],y[2]);
    CSA     CSA_240_336(c2[3],ip2[2],ip1[3],c1[3],x[3],y[2]);
    CSA     CSA_320_336(c2[4],ip2[3],ip1[4],c1[4],x[4],y[2]);
    CSA     CSA_400_336(c2[5],ip2[4],ip1[5],c1[5],x[5],y[2]);
    CSA     CSA_480_336(c2[6],ip2[5],ip1[6],c1[6],x[6],y[2]);
    CSA     CSA_560_336(c2[7],ip2[6],ip1[7],c1[7],x[7],y[2]);
    CSA     CSA_640_336(c2[8],ip2[7],ip1[8],c1[8],x[8],y[2]);
    CSA     CSA_720_336(c2[9],ip2[8],ip1[9],c1[9],x[9],y[2]);
    CSA     CSA_800_336(c2[10],ip2[9],ip1[10],c1[10],x[10],y[2]);
    CSA     CSA_880_336(c2[11],ip2[10],ip1[11],c1[11],x[11],y[2]);
    CSA     CSA_960_336(c2[12],ip2[11],ip1[12],c1[12],x[12],y[2]);
    CSA     CSA_1040_336(c2[13],ip2[12],ip1[13],c1[13],x[13],y[2]);
    CSA     CSA_1120_336(c2[14],ip2[13],ip1[14],c1[14],x[14],y[2]);
    CSA     CSA_1200_336(c2[15],ip2[14],1'b0  ,c1[15],x[15],y[2]);
    CSA     CSA_0_504(c3[0],p  [3],ip2[0],c2[0],x[0],y[3]);
    CSA     CSA_80_504(c3[1],ip3[0],ip2[1],c2[1],x[1],y[3]);
    CSA     CSA_160_504(c3[2],ip3[1],ip2[2],c2[2],x[2],y[3]);
    CSA     CSA_240_504(c3[3],ip3[2],ip2[3],c2[3],x[3],y[3]);
    CSA     CSA_320_504(c3[4],ip3[3],ip2[4],c2[4],x[4],y[3]);
    CSA     CSA_400_504(c3[5],ip3[4],ip2[5],c2[5],x[5],y[3]);
    CSA     CSA_480_504(c3[6],ip3[5],ip2[6],c2[6],x[6],y[3]);
    CSA     CSA_560_504(c3[7],ip3[6],ip2[7],c2[7],x[7],y[3]);
    CSA     CSA_640_504(c3[8],ip3[7],ip2[8],c2[8],x[8],y[3]);
    CSA     CSA_720_504(c3[9],ip3[8],ip2[9],c2[9],x[9],y[3]);
    CSA     CSA_800_504(c3[10],ip3[9],ip2[10],c2[10],x[10],y[3]);
    CSA     CSA_880_504(c3[11],ip3[10],ip2[11],c2[11],x[11],y[3]);
    CSA     CSA_960_504(c3[12],ip3[11],ip2[12],c2[12],x[12],y[3]);
    CSA     CSA_1040_504(c3[13],ip3[12],ip2[13],c2[13],x[13],y[3]);
    CSA     CSA_1120_504(c3[14],ip3[13],ip2[14],c2[14],x[14],y[3]);
    CSA     CSA_1200_504(c3[15],ip3[14],1'b0  ,c2[15],x[15],y[3]);
    CSA     CSA_0_672(c4[0],p  [4],ip3[0],c3[0],x[0],y[4]);
    CSA     CSA_80_672(c4[1],ip4[0],ip3[1],c3[1],x[1],y[4]);
    CSA     CSA_160_672(c4[2],ip4[1],ip3[2],c3[2],x[2],y[4]);
    CSA     CSA_240_672(c4[3],ip4[2],ip3[3],c3[3],x[3],y[4]);
    CSA     CSA_320_672(c4[4],ip4[3],ip3[4],c3[4],x[4],y[4]);
    CSA     CSA_400_672(c4[5],ip4[4],ip3[5],c3[5],x[5],y[4]);
    CSA     CSA_480_672(c4[6],ip4[5],ip3[6],c3[6],x[6],y[4]);
    CSA     CSA_560_672(c4[7],ip4[6],ip3[7],c3[7],x[7],y[4]);
    CSA     CSA_640_672(c4[8],ip4[7],ip3[8],c3[8],x[8],y[4]);
    CSA     CSA_720_672(c4[9],ip4[8],ip3[9],c3[9],x[9],y[4]);
    CSA     CSA_800_672(c4[10],ip4[9],ip3[10],c3[10],x[10],y[4]);
    CSA     CSA_880_672(c4[11],ip4[10],ip3[11],c3[11],x[11],y[4]);
    CSA     CSA_960_672(c4[12],ip4[11],ip3[12],c3[12],x[12],y[4]);
    CSA     CSA_1040_672(c4[13],ip4[12],ip3[13],c3[13],x[13],y[4]);
    CSA     CSA_1120_672(c4[14],ip4[13],ip3[14],c3[14],x[14],y[4]);
    CSA     CSA_1200_672(c4[15],ip4[14],1'b0  ,c3[15],x[15],y[4]);
    CSA     CSA_0_840(c5[0],p  [5],ip4[0],c4[0],x[0],y[5]);
    CSA     CSA_80_840(c5[1],ip5[0],ip4[1],c4[1],x[1],y[5]);
    CSA     CSA_160_840(c5[2],ip5[1],ip4[2],c4[2],x[2],y[5]);
    CSA     CSA_240_840(c5[3],ip5[2],ip4[3],c4[3],x[3],y[5]);
    CSA     CSA_320_840(c5[4],ip5[3],ip4[4],c4[4],x[4],y[5]);
    CSA     CSA_400_840(c5[5],ip5[4],ip4[5],c4[5],x[5],y[5]);
    CSA     CSA_480_840(c5[6],ip5[5],ip4[6],c4[6],x[6],y[5]);
    CSA     CSA_560_840(c5[7],ip5[6],ip4[7],c4[7],x[7],y[5]);
    CSA     CSA_640_840(c5[8],ip5[7],ip4[8],c4[8],x[8],y[5]);
    CSA     CSA_720_840(c5[9],ip5[8],ip4[9],c4[9],x[9],y[5]);
    CSA     CSA_800_840(c5[10],ip5[9],ip4[10],c4[10],x[10],y[5]);
    CSA     CSA_880_840(c5[11],ip5[10],ip4[11],c4[11],x[11],y[5]);
    CSA     CSA_960_840(c5[12],ip5[11],ip4[12],c4[12],x[12],y[5]);
    CSA     CSA_1040_840(c5[13],ip5[12],ip4[13],c4[13],x[13],y[5]);
    CSA     CSA_1120_840(c5[14],ip5[13],ip4[14],c4[14],x[14],y[5]);
    CSA     CSA_1200_840(c5[15],ip5[14],1'b0  ,c4[15],x[15],y[5]);
    CSA     CSA_0_1008(c6[0],p  [6],ip5[0],c5[0],x[0],y[6]);
    CSA     CSA_80_1008(c6[1],ip6[0],ip5[1],c5[1],x[1],y[6]);
    CSA     CSA_160_1008(c6[2],ip6[1],ip5[2],c5[2],x[2],y[6]);
    CSA     CSA_240_1008(c6[3],ip6[2],ip5[3],c5[3],x[3],y[6]);
    CSA     CSA_320_1008(c6[4],ip6[3],ip5[4],c5[4],x[4],y[6]);
    CSA     CSA_400_1008(c6[5],ip6[4],ip5[5],c5[5],x[5],y[6]);
    CSA     CSA_480_1008(c6[6],ip6[5],ip5[6],c5[6],x[6],y[6]);
    CSA     CSA_560_1008(c6[7],ip6[6],ip5[7],c5[7],x[7],y[6]);
    CSA     CSA_640_1008(c6[8],ip6[7],ip5[8],c5[8],x[8],y[6]);
    CSA     CSA_720_1008(c6[9],ip6[8],ip5[9],c5[9],x[9],y[6]);
    CSA     CSA_800_1008(c6[10],ip6[9],ip5[10],c5[10],x[10],y[6]);
    CSA     CSA_880_1008(c6[11],ip6[10],ip5[11],c5[11],x[11],y[6]);
    CSA     CSA_960_1008(c6[12],ip6[11],ip5[12],c5[12],x[12],y[6]);
    CSA     CSA_1040_1008(c6[13],ip6[12],ip5[13],c5[13],x[13],y[6]);
    CSA     CSA_1120_1008(c6[14],ip6[13],ip5[14],c5[14],x[14],y[6]);
    CSA     CSA_1200_1008(c6[15],ip6[14],1'b0  ,c5[15],x[15],y[6]);
    CSA     CSA_0_1176(c7[0],p  [7],ip6[0],c6[0],x[0],y[7]);
    CSA     CSA_80_1176(c7[1],ip7[0],ip6[1],c6[1],x[1],y[7]);
    CSA     CSA_160_1176(c7[2],ip7[1],ip6[2],c6[2],x[2],y[7]);
    CSA     CSA_240_1176(c7[3],ip7[2],ip6[3],c6[3],x[3],y[7]);
    CSA     CSA_320_1176(c7[4],ip7[3],ip6[4],c6[4],x[4],y[7]);
    CSA     CSA_400_1176(c7[5],ip7[4],ip6[5],c6[5],x[5],y[7]);
    CSA     CSA_480_1176(c7[6],ip7[5],ip6[6],c6[6],x[6],y[7]);
    CSA     CSA_560_1176(c7[7],ip7[6],ip6[7],c6[7],x[7],y[7]);
    CSA     CSA_640_1176(c7[8],ip7[7],ip6[8],c6[8],x[8],y[7]);
    CSA     CSA_720_1176(c7[9],ip7[8],ip6[9],c6[9],x[9],y[7]);
    CSA     CSA_800_1176(c7[10],ip7[9],ip6[10],c6[10],x[10],y[7]);
    CSA     CSA_880_1176(c7[11],ip7[10],ip6[11],c6[11],x[11],y[7]);
    CSA     CSA_960_1176(c7[12],ip7[11],ip6[12],c6[12],x[12],y[7]);
    CSA     CSA_1040_1176(c7[13],ip7[12],ip6[13],c6[13],x[13],y[7]);
    CSA     CSA_1120_1176(c7[14],ip7[13],ip6[14],c6[14],x[14],y[7]);
    CSA     CSA_1200_1176(c7[15],ip7[14],1'b0  ,c6[15],x[15],y[7]);
    CSA     CSA_0_1344(c8[0],p  [8],ip7[0],c7[0],x[0],y[8]);
    CSA     CSA_80_1344(c8[1],ip8[0],ip7[1],c7[1],x[1],y[8]);
    CSA     CSA_160_1344(c8[2],ip8[1],ip7[2],c7[2],x[2],y[8]);
    CSA     CSA_240_1344(c8[3],ip8[2],ip7[3],c7[3],x[3],y[8]);
    CSA     CSA_320_1344(c8[4],ip8[3],ip7[4],c7[4],x[4],y[8]);
    CSA     CSA_400_1344(c8[5],ip8[4],ip7[5],c7[5],x[5],y[8]);
    CSA     CSA_480_1344(c8[6],ip8[5],ip7[6],c7[6],x[6],y[8]);
    CSA     CSA_560_1344(c8[7],ip8[6],ip7[7],c7[7],x[7],y[8]);
    CSA     CSA_640_1344(c8[8],ip8[7],ip7[8],c7[8],x[8],y[8]);
    CSA     CSA_720_1344(c8[9],ip8[8],ip7[9],c7[9],x[9],y[8]);
    CSA     CSA_800_1344(c8[10],ip8[9],ip7[10],c7[10],x[10],y[8]);
    CSA     CSA_880_1344(c8[11],ip8[10],ip7[11],c7[11],x[11],y[8]);
    CSA     CSA_960_1344(c8[12],ip8[11],ip7[12],c7[12],x[12],y[8]);
    CSA     CSA_1040_1344(c8[13],ip8[12],ip7[13],c7[13],x[13],y[8]);
    CSA     CSA_1120_1344(c8[14],ip8[13],ip7[14],c7[14],x[14],y[8]);
    CSA     CSA_1200_1344(c8[15],ip8[14],1'b0  ,c7[15],x[15],y[8]);
    CSA     CSA_0_1512(c9[0],p  [9],ip8[0],c8[0],x[0],y[9]);
    CSA     CSA_80_1512(c9[1],ip9[0],ip8[1],c8[1],x[1],y[9]);
    CSA     CSA_160_1512(c9[2],ip9[1],ip8[2],c8[2],x[2],y[9]);
    CSA     CSA_240_1512(c9[3],ip9[2],ip8[3],c8[3],x[3],y[9]);
    CSA     CSA_320_1512(c9[4],ip9[3],ip8[4],c8[4],x[4],y[9]);
    CSA     CSA_400_1512(c9[5],ip9[4],ip8[5],c8[5],x[5],y[9]);
    CSA     CSA_480_1512(c9[6],ip9[5],ip8[6],c8[6],x[6],y[9]);
    CSA     CSA_560_1512(c9[7],ip9[6],ip8[7],c8[7],x[7],y[9]);
    CSA     CSA_640_1512(c9[8],ip9[7],ip8[8],c8[8],x[8],y[9]);
    CSA     CSA_720_1512(c9[9],ip9[8],ip8[9],c8[9],x[9],y[9]);
    CSA     CSA_800_1512(c9[10],ip9[9],ip8[10],c8[10],x[10],y[9]);
    CSA     CSA_880_1512(c9[11],ip9[10],ip8[11],c8[11],x[11],y[9]);
    CSA     CSA_960_1512(c9[12],ip9[11],ip8[12],c8[12],x[12],y[9]);
    CSA     CSA_1040_1512(c9[13],ip9[12],ip8[13],c8[13],x[13],y[9]);
    CSA     CSA_1120_1512(c9[14],ip9[13],ip8[14],c8[14],x[14],y[9]);
    CSA     CSA_1200_1512(c9[15],ip9[14],1'b0  ,c8[15],x[15],y[9]);
    CSA     CSA_0_1680(c10[0],p  [10],ip9[0],c9[0],x[0],y[10]);
    CSA     CSA_80_1680(c10[1],ip10[0],ip9[1],c9[1],x[1],y[10]);
    CSA     CSA_160_1680(c10[2],ip10[1],ip9[2],c9[2],x[2],y[10]);
    CSA     CSA_240_1680(c10[3],ip10[2],ip9[3],c9[3],x[3],y[10]);
    CSA     CSA_320_1680(c10[4],ip10[3],ip9[4],c9[4],x[4],y[10]);
    CSA     CSA_400_1680(c10[5],ip10[4],ip9[5],c9[5],x[5],y[10]);
    CSA     CSA_480_1680(c10[6],ip10[5],ip9[6],c9[6],x[6],y[10]);
    CSA     CSA_560_1680(c10[7],ip10[6],ip9[7],c9[7],x[7],y[10]);
    CSA     CSA_640_1680(c10[8],ip10[7],ip9[8],c9[8],x[8],y[10]);
    CSA     CSA_720_1680(c10[9],ip10[8],ip9[9],c9[9],x[9],y[10]);
    CSA     CSA_800_1680(c10[10],ip10[9],ip9[10],c9[10],x[10],y[10]);
    CSA     CSA_880_1680(c10[11],ip10[10],ip9[11],c9[11],x[11],y[10]);
    CSA     CSA_960_1680(c10[12],ip10[11],ip9[12],c9[12],x[12],y[10]);
    CSA     CSA_1040_1680(c10[13],ip10[12],ip9[13],c9[13],x[13],y[10]);
    CSA     CSA_1120_1680(c10[14],ip10[13],ip9[14],c9[14],x[14],y[10]);
    CSA     CSA_1200_1680(c10[15],ip10[14],1'b0  ,c9[15],x[15],y[10]);
    CSA     CSA_0_1848(c11[0],p  [11],ip10[0],c10[0],x[0],y[11]);
    CSA     CSA_80_1848(c11[1],ip11[0],ip10[1],c10[1],x[1],y[11]);
    CSA     CSA_160_1848(c11[2],ip11[1],ip10[2],c10[2],x[2],y[11]);
    CSA     CSA_240_1848(c11[3],ip11[2],ip10[3],c10[3],x[3],y[11]);
    CSA     CSA_320_1848(c11[4],ip11[3],ip10[4],c10[4],x[4],y[11]);
    CSA     CSA_400_1848(c11[5],ip11[4],ip10[5],c10[5],x[5],y[11]);
    CSA     CSA_480_1848(c11[6],ip11[5],ip10[6],c10[6],x[6],y[11]);
    CSA     CSA_560_1848(c11[7],ip11[6],ip10[7],c10[7],x[7],y[11]);
    CSA     CSA_640_1848(c11[8],ip11[7],ip10[8],c10[8],x[8],y[11]);
    CSA     CSA_720_1848(c11[9],ip11[8],ip10[9],c10[9],x[9],y[11]);
    CSA     CSA_800_1848(c11[10],ip11[9],ip10[10],c10[10],x[10],y[11]);
    CSA     CSA_880_1848(c11[11],ip11[10],ip10[11],c10[11],x[11],y[11]);
    CSA     CSA_960_1848(c11[12],ip11[11],ip10[12],c10[12],x[12],y[11]);
    CSA     CSA_1040_1848(c11[13],ip11[12],ip10[13],c10[13],x[13],y[11]);
    CSA     CSA_1120_1848(c11[14],ip11[13],ip10[14],c10[14],x[14],y[11]);
    CSA     CSA_1200_1848(c11[15],ip11[14],1'b0  ,c10[15],x[15],y[11]);
    CSA     CSA_0_2016(c12[0],p  [12],ip11[0],c11[0],x[0],y[12]);
    CSA     CSA_80_2016(c12[1],ip12[0],ip11[1],c11[1],x[1],y[12]);
    CSA     CSA_160_2016(c12[2],ip12[1],ip11[2],c11[2],x[2],y[12]);
    CSA     CSA_240_2016(c12[3],ip12[2],ip11[3],c11[3],x[3],y[12]);
    CSA     CSA_320_2016(c12[4],ip12[3],ip11[4],c11[4],x[4],y[12]);
    CSA     CSA_400_2016(c12[5],ip12[4],ip11[5],c11[5],x[5],y[12]);
    CSA     CSA_480_2016(c12[6],ip12[5],ip11[6],c11[6],x[6],y[12]);
    CSA     CSA_560_2016(c12[7],ip12[6],ip11[7],c11[7],x[7],y[12]);
    CSA     CSA_640_2016(c12[8],ip12[7],ip11[8],c11[8],x[8],y[12]);
    CSA     CSA_720_2016(c12[9],ip12[8],ip11[9],c11[9],x[9],y[12]);
    CSA     CSA_800_2016(c12[10],ip12[9],ip11[10],c11[10],x[10],y[12]);
    CSA     CSA_880_2016(c12[11],ip12[10],ip11[11],c11[11],x[11],y[12]);
    CSA     CSA_960_2016(c12[12],ip12[11],ip11[12],c11[12],x[12],y[12]);
    CSA     CSA_1040_2016(c12[13],ip12[12],ip11[13],c11[13],x[13],y[12]);
    CSA     CSA_1120_2016(c12[14],ip12[13],ip11[14],c11[14],x[14],y[12]);
    CSA     CSA_1200_2016(c12[15],ip12[14],1'b0  ,c11[15],x[15],y[12]);
    CSA     CSA_0_2184(c13[0],p  [13],ip12[0],c12[0],x[0],y[13]);
    CSA     CSA_80_2184(c13[1],ip13[0],ip12[1],c12[1],x[1],y[13]);
    CSA     CSA_160_2184(c13[2],ip13[1],ip12[2],c12[2],x[2],y[13]);
    CSA     CSA_240_2184(c13[3],ip13[2],ip12[3],c12[3],x[3],y[13]);
    CSA     CSA_320_2184(c13[4],ip13[3],ip12[4],c12[4],x[4],y[13]);
    CSA     CSA_400_2184(c13[5],ip13[4],ip12[5],c12[5],x[5],y[13]);
    CSA     CSA_480_2184(c13[6],ip13[5],ip12[6],c12[6],x[6],y[13]);
    CSA     CSA_560_2184(c13[7],ip13[6],ip12[7],c12[7],x[7],y[13]);
    CSA     CSA_640_2184(c13[8],ip13[7],ip12[8],c12[8],x[8],y[13]);
    CSA     CSA_720_2184(c13[9],ip13[8],ip12[9],c12[9],x[9],y[13]);
    CSA     CSA_800_2184(c13[10],ip13[9],ip12[10],c12[10],x[10],y[13]);
    CSA     CSA_880_2184(c13[11],ip13[10],ip12[11],c12[11],x[11],y[13]);
    CSA     CSA_960_2184(c13[12],ip13[11],ip12[12],c12[12],x[12],y[13]);
    CSA     CSA_1040_2184(c13[13],ip13[12],ip12[13],c12[13],x[13],y[13]);
    CSA     CSA_1120_2184(c13[14],ip13[13],ip12[14],c12[14],x[14],y[13]);
    CSA     CSA_1200_2184(c13[15],ip13[14],1'b0  ,c12[15],x[15],y[13]);
    CSA     CSA_0_2352(c14[0],p  [14],ip13[0],c13[0],x[0],y[14]);
    CSA     CSA_80_2352(c14[1],ip14[0],ip13[1],c13[1],x[1],y[14]);
    CSA     CSA_160_2352(c14[2],ip14[1],ip13[2],c13[2],x[2],y[14]);
    CSA     CSA_240_2352(c14[3],ip14[2],ip13[3],c13[3],x[3],y[14]);
    CSA     CSA_320_2352(c14[4],ip14[3],ip13[4],c13[4],x[4],y[14]);
    CSA     CSA_400_2352(c14[5],ip14[4],ip13[5],c13[5],x[5],y[14]);
    CSA     CSA_480_2352(c14[6],ip14[5],ip13[6],c13[6],x[6],y[14]);
    CSA     CSA_560_2352(c14[7],ip14[6],ip13[7],c13[7],x[7],y[14]);
    CSA     CSA_640_2352(c14[8],ip14[7],ip13[8],c13[8],x[8],y[14]);
    CSA     CSA_720_2352(c14[9],ip14[8],ip13[9],c13[9],x[9],y[14]);
    CSA     CSA_800_2352(c14[10],ip14[9],ip13[10],c13[10],x[10],y[14]);
    CSA     CSA_880_2352(c14[11],ip14[10],ip13[11],c13[11],x[11],y[14]);
    CSA     CSA_960_2352(c14[12],ip14[11],ip13[12],c13[12],x[12],y[14]);
    CSA     CSA_1040_2352(c14[13],ip14[12],ip13[13],c13[13],x[13],y[14]);
    CSA     CSA_1120_2352(c14[14],ip14[13],ip13[14],c13[14],x[14],y[14]);
    CSA     CSA_1200_2352(c14[15],ip14[14],1'b0  ,c13[15],x[15],y[14]);
    CSA     CSA_0_2520(c15[0],p  [15],ip14[0],c14[0],x[0],y[15]);
    CSA     CSA_80_2520(c15[1],ip15[0],ip14[1],c14[1],x[1],y[15]);
    CSA     CSA_160_2520(c15[2],ip15[1],ip14[2],c14[2],x[2],y[15]);
    CSA     CSA_240_2520(c15[3],ip15[2],ip14[3],c14[3],x[3],y[15]);
    CSA     CSA_320_2520(c15[4],ip15[3],ip14[4],c14[4],x[4],y[15]);
    CSA     CSA_400_2520(c15[5],ip15[4],ip14[5],c14[5],x[5],y[15]);
    CSA     CSA_480_2520(c15[6],ip15[5],ip14[6],c14[6],x[6],y[15]);
    CSA     CSA_560_2520(c15[7],ip15[6],ip14[7],c14[7],x[7],y[15]);
    CSA     CSA_640_2520(c15[8],ip15[7],ip14[8],c14[8],x[8],y[15]);
    CSA     CSA_720_2520(c15[9],ip15[8],ip14[9],c14[9],x[9],y[15]);
    CSA     CSA_800_2520(c15[10],ip15[9],ip14[10],c14[10],x[10],y[15]);
    CSA     CSA_880_2520(c15[11],ip15[10],ip14[11],c14[11],x[11],y[15]);
    CSA     CSA_960_2520(c15[12],ip15[11],ip14[12],c14[12],x[12],y[15]);
    CSA     CSA_1040_2520(c15[13],ip15[12],ip14[13],c14[13],x[13],y[15]);
    CSA     CSA_1120_2520(c15[14],ip15[13],ip14[14],c14[14],x[14],y[15]);
    CSA     CSA_1200_2520(c15[15],ip15[14],1'b0  ,c14[15],x[15],y[15]);
    fullAdd FA_0_2688(c16[0],p[16],ip15[0],c15[0],1'b0 );
    fullAdd FA_80_2688(c16[1],p[17],ip15[1],c15[1],c16[0]);
    fullAdd FA_160_2688(c16[2],p[18],ip15[2],c15[2],c16[1]);
    fullAdd FA_240_2688(c16[3],p[19],ip15[3],c15[3],c16[2]);
    fullAdd FA_320_2688(c16[4],p[20],ip15[4],c15[4],c16[3]);
    fullAdd FA_400_2688(c16[5],p[21],ip15[5],c15[5],c16[4]);
    fullAdd FA_480_2688(c16[6],p[22],ip15[6],c15[6],c16[5]);
    fullAdd FA_560_2688(c16[7],p[23],ip15[7],c15[7],c16[6]);
    fullAdd FA_640_2688(c16[8],p[24],ip15[8],c15[8],c16[7]);
    fullAdd FA_720_2688(c16[9],p[25],ip15[9],c15[9],c16[8]);
    fullAdd FA_800_2688(c16[10],p[26],ip15[10],c15[10],c16[9]);
    fullAdd FA_880_2688(c16[11],p[27],ip15[11],c15[11],c16[10]);
    fullAdd FA_960_2688(c16[12],p[28],ip15[12],c15[12],c16[11]);
    fullAdd FA_1040_2688(c16[13],p[29],ip15[13],c15[13],c16[12]);
    fullAdd FA_1120_2688(c16[14],p[30],ip15[14],c15[14],c16[13]);
    fullAdd FA_1200_2688(c16[15],p[31],1'b0  ,c15[15],c16[14]);
endmodule
